-- LCS-2016-099: Extended Ranges
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_099
-- TODO
