-- LCS-2016-050: API for Assert
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_050
-- TODO
