-- LCS-2016-030: Garbage Collection
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_030
-- TODO
