-- LCS-2016-026c: Long Integers
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_026c

package pack026c is

    constant a : integer := 89345897098345;
    constant b : integer := -892348978489894 ;

    constant c : natural := 723478927649492389 ;

end package;
