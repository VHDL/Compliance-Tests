-- LCS-2016-082: Empty Record
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_082

package pack is

    record rec is
    end record ;

end package;
