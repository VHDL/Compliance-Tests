-- LCS-2016-082: Empty Record
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_082

package pack082 is

    type rec is record
    end record ;

end package;
