-- LCS-2016-034: Attributes for PSL
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_043
-- TODO
