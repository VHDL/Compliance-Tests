-- LCS-2016-071a: Extra optional semicolon at the end of interface_list
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_071a
entity e071a is
  port (
    a   :   in  bit ;
    b   :   out integer ;
  ) ;
end entity ;

--

library vunit_lib;
context vunit_lib.vunit_context;

entity tb_extra_optional_semicolon_on_interface_list is
  generic ( runner_cfg : string );
end entity;

architecture tb of tb_extra_optional_semicolon_on_interface_list is
begin
  test_runner: process is
  begin
    test_runner_setup(runner, runner_cfg);
    info("LCS-2016-071a: Extra optional semicolon at the end of interface list");
    test_runner_cleanup(runner);
    wait;
  end process test_runner;
end architecture tb;
