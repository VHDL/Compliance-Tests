-- LCS-2016-045c: Interface - 'CONVERSE for a mode view
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_045c
-- TODO
