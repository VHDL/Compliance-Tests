-- LCS-2016-011: Date/Time Functions
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_011
-- TODO
