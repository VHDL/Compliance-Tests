-- LCS-2016-061: Conditional Compilation
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_061
-- TODO
