-- LCS-2016-018: Attributes for Enumerated Types
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_018
-- TODO
