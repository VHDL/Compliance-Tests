-- LCS-2016-072b: Function knows return vector size
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_072b
-- TODO
