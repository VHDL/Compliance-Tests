context vunit_context is
  library vunit_lib;
  use vunit_lib.mock_pkg.all;
  use vunit_lib.check_equal_pkg.all;
end context;
