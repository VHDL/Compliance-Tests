-- LCS-2016-002: Allow access and protected type parameters on function interfaces
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_002
-- TODO
