-- LCS-2016-018d: New attribute - 'DESGINATED_TYPE
-- http://www.eda-twiki.org/cgi-bin/view.cgi/P1076/LCS2016_018d
-- TODO
